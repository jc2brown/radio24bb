`timescale 1ps / 1ps

module tb_fir_filter(

    );
    
    

    
        
wire [31:0] sig_p;
    
siggen
#(
    .AMPL(127e-6),
    .FREQ(1e7)
)
siggen_a 
(
    .sig_p_uv(sig_p)
);
    
    
    
    
    
reg clk = 1'b1;
always #5000 clk <= !clk;

reg reset = 1'b1;
initial #100000 reset <= 1'b0;
    

reg [1:0] valid_in = 2'h3;
//always @(posedge clk) valid_in <= valid_in + 1;

wire [7:0] out;
wire valid_out;


reg [24:0] cfg_din = 'h0;
reg cfg_ce = 1'b0;
    
wire [17:0] in = sig_p;
//wire [17:0] in = { {11{!sig_p[7]}}, {7{sig_p[7]}} };

fir_filter #( .LEN(21) ) 
dut (    
    .reset(reset),
    .clk(clk),

    .cfg_din(cfg_din),
    .cfg_ce(cfg_ce),
    
    .len(),    

    .in(&valid_in ? in : 0),
    .valid_in(&valid_in),
    
    .out(out),
    .valid_out(valid_out)

);
    
    
    
real coef[0:20] = {    
/*
    0.018121627, -0.0025737102, -0.049848193,
	-0.048790703, 0.046189787, 0.086422509, -0.075657994, -0.24352923, -0.050645060,
	0.45368918, 0.73324356, 0.45368918, -0.050645060, -0.24352923, -0.075657994,
	0.086422509, 0.046189787, -0.048790703, -0.049848193, -0.0025737102, 0.018121627
	*/
	/*
	0.0020676081, -0.0010862434, -0.028109706,
        -0.015849916, 0.0067964367, 0.0043629139, 0.015229101, -0.12102499, -0.24878713,
        0.37998359, 1.0128367, 0.37998359, -0.24878713, -0.12102499, 0.015229101,
        0.0043629139, 0.0067964367, -0.015849916, -0.028109706, -0.0010862434, 0.0020676081
        */
        /*
      0.000019538157, 0.000029681056, 0.000016285841,
            0.000045572917, 0.000013777408, 0.000085082212, 0.000012272895, 0.00022904898, 0.000011470952,
            0.0020298291, 0.99501488, 0.0020298291, 0.000011470952, 0.00022904898, 0.000012272895,
            0.000085082212, 0.000013777408, 0.000045572917, 0.000016285841, 0.000029681056, 0.000019538157,
            */
            
            
            1.1, 
            0.0, 0.0, 0.0, 0.0, 0.0, 
            0.0, 0.0, 0.0, 0.0, 0.0, 
            0.0, 0.0, 0.0, 0.0, 0.0,
            0.0, 0.0, 0.0, 0.0, 0.0
            
};
	
	
	
reg [7:0] x;
always @(posedge clk) if (valid_out) x <= out;

	
integer i;    
    
initial begin

    @(negedge reset);

    @(posedge clk) begin
        cfg_din <= $rtoi(2**23 * coef[0]);
        cfg_ce <= 1;
    end
    
    
    for (i=1; i<21; i=i+1) begin
        @(posedge clk) cfg_din <= $rtoi(2**23 * coef[i]);
    end
    
    
    @(posedge clk) cfg_ce <= 1'b0;
/*
	0.052575624, 1.9468305, 0.052575624, -0.050807312, 0.047904049, -0.043930688,
	0.038975989, -0.033150630, 0.026584741, -0.019424993, 0.011831323, -0.0039733604
*/



end
    
    
    
    
    
endmodule

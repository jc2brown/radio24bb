
/*


package tb_utils;
    
    
        
         
        
endpackage


*/